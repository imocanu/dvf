package dvf_lib_pkg;
  import uvm_pkg::*;

  `include "uvm_macros.svh"

  string msg_id = "dvf_lib";

  `include "dvf_agent_cfg.sv"
  `include "dvf_monitor.sv"
  `include "dvf_sequencer.sv"
  `include "dvf_driver.sv"
  `include "dvf_agent.sv"
  `include "dvf_seq.sv"
  `include "dvf_env_cfg.sv"
  `include "dvf_virtual_sequencer.sv"
  `include "dvf_scoreboard.sv"
  `include "dvf_env.sv"
  `include "dvf_vseq.sv"
  `include "dvf_test.sv"

endpackage